module hello_world();
initial begin
$display("\n Hello angel\n");
end
endmodule