module helloworld();
  initial begin
    $display("\n Hello World! \n");
  end
endmodule
